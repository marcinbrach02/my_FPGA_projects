module tester_module(







);
endmodule
 