module microSD(
	input wire clk,
	input wire rst,
	input wire cs,
	input wire [47:0] command 
	
);


//case do obs�ugi rozkazu do karty poprzez wys�anie komendy?






endmodule